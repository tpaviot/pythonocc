--  Copyright (C) 2007-2008  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--
-- File:	GEOMAlgo_Tools3D.cdl
-- Created:	
-- Author:	Peter KURNEV  
--
class Tools3D from GEOMAlgo 

	---Purpose:  Auxiliary tools for Algorithms   

uses  
    State     from TopAbs,
    ShapeEnum from TopAbs, 
    Pnt from gp, 
    Shape  from TopoDS, 
    Vertex from TopoDS,
    Edge   from TopoDS, 
    Face   from TopoDS,  
    Solid  from TopoDS, 
     
    ListOfShape       from TopTools, 
    IndexedMapOfShape from TopTools, 
    IndexedDataMapOfShapeListOfShape from TopTools, 
    Context from IntTools,  
    ListOfCoupleOfShape from NMTTools
    
--raises

is 
    IsSplitToReverse(myclass;  
		theSplit   :  Shape from TopoDS; 
		theShape   :  Shape from TopoDS; 
    	    	theContext:out Context from IntTools)  
    	---Purpose: Returns True if the shape theSplit has opposite 
    	--          direction than theShape 
	--          theContext - cashed geometrical tools
    	returns Boolean from Standard; 
	 
    IsSplitToReverse(myclass;  
		theSplit  :  Face from TopoDS; 
		theShape  :  Face from TopoDS; 
    	    	theContext:out Context from IntTools) 
    	---Purpose: Returns True if normal direction of the face   
    	--          theShape is not the same as for the face  
    	--          theSplit 
        --          theContext - cashed geometrical tools 
    	returns Boolean from Standard; 
     
    IsSplitToReverse(myclass;  
		theEdge   :  Edge from TopoDS; 
		theSplit  :  Edge from TopoDS; 
    	    	theContext:out Context from IntTools) 
    	---Purpose: Returns True if tangent direction of the edge   
    	--          theEdge is not the same as for the edge  
    	--          theSplit    
	--          theContext - cashed geometrical tools 
    	returns Boolean from Standard;  
	 
    Sense  (myclass;  
    	    	theF1:  Face from TopoDS; 
	    	theF2:  Face from TopoDS) 
	---Purpose: For the couple of faces theF1, theF2 
	--          computes sense value      		 
	--          Returns 0 if the faces are not sensible         		 
	--          Returns 1 if the faces have same sense         		 
	--          Returns 2 if the faces have opposite sense         		 
	returns Integer from Standard; 

    CopyFace(myclass;  
    	    	theF1:  Face from TopoDS; 
	    	theF2:out Face from TopoDS); 
    	---Purpose: Makes new face theF2 from surface and wires  
    	--          of the face theF1 
	 
    MakeContainer(myclass; 
    	    	theType:ShapeEnum from TopAbs; 
		theShape:out Shape from TopoDS); 
	---Purpose: Makes empty shape theShape of the type theType        
		 
		
    MakeConnexityBlock(myclass; 
                theLS      :ListOfShape from TopTools;   
		theMapAvoid:IndexedMapOfShape from TopTools;       		 
		theLSCB    :out ListOfShape from TopTools);   
    	---Purpose: For the list of faces theLS build block  
    	--          theLSCB in terms of connexity by edges   
        --          theMapAvoid - set of edges to avoid for 
	--          the treatment 
	
    ComputeStateByOnePoint(myclass; 
    	    	theShape :Shape from TopoDS;  
    	    	theSolid :Solid from TopoDS;  
		theTol   :Real from Standard;       
    	    	theContext:out Context from IntTools) 
    	---Purpose: Computes the 3-D state of the shape theShape 
	--          toward solid theSolid. 
	--          theTol - value of precision of computation   
        --          theContext- cahed geometrical tools  
        --          Returns 3-D state. 
    	returns State from TopAbs;  

    ComputeState(myclass; 
    	    	thePoint :Pnt  from gp;  
    	    	theSolid :Solid from TopoDS;  
		theTol   :Real from Standard;       
    	    	theContext:out Context from IntTools) 
	---Purpose: Computes the 3-D state of the point thePoint 
	--          toward solid theSolid. 
	--          theTol - value of precision of computation   
        --          theContext- cahed geometrical tools  
        --          Returns 3-D state. 
     	returns State from TopAbs;  
	
    ComputeState(myclass; 
    	    	theVertex:Vertex from TopoDS;  
    	    	theSolid :Solid from TopoDS;  
		theTol   :Real from Standard;       
    	    	theContext:out Context from IntTools) 
    	---Purpose: Computes the 3-D state of the vertex theVertex 
	--          toward solid theSolid. 
	--          theTol - value of precision of computation   
        --          theContext- cahed geometrical tools  
        --          Returns 3-D state. 
	returns State from TopAbs;  
	
    ComputeState(myclass; 
    	    	theEdge  :Edge  from TopoDS;  
    	    	theSolid :Solid from TopoDS;  
		theTol   :Real from Standard;       
    	    	theContext:out Context from IntTools) 
	---Purpose: Computes the 3-D state of the edge theEdge 
	--          toward solid theSolid. 
	--          theTol - value of precision of computation   
        --          theContext- cahed geometrical tools  
        --          Returns 3-D state. 
	returns State from TopAbs;  
	
    ComputeState(myclass; 
    	    	theFace  :Face  from TopoDS;  
    	    	theSolid :Solid from TopoDS;  
		theTol   :Real from Standard;  
                theBounds:IndexedMapOfShape from TopTools; 		 
    	    	theContext:out Context from IntTools) 
    	---Purpose: Computes the 3-D state of the face theFace 
	--          toward solid theSolid. 
	--          theTol - value of precision of computation   
        --          theBounds - set of edges of theFace to avoid          
        --          theContext- cahed geometrical tools  
        --          Returns 3-D state. 
    	returns State from TopAbs; 

    IsInternalFace(myclass; 
    	    	theFace  :Face from TopoDS; 
    	    	theEdge  :Edge from TopoDS; 
    	    	theFace1 :Face from TopoDS; 
    	    	theFace2 :Face from TopoDS) 
    	---Purpose: Returns True if the face theFace is inside of the  
	--          couple of faces theFace1, theFace2. 
	--          The faces theFace, theFace1, theFace2  must 
        --          share the edge theEdge  	 
    	returns Boolean from Standard; 
	 
    IsInternalFace(myclass; 
    	    	theFace :Face  from TopoDS; 
    	    	theEdge :Edge  from TopoDS; 
    	    	theLF   :ListOfShape from TopTools)  
    	---Purpose: Returns True if the face theFace is inside of the  
	--          appropriate couple of faces (from the set theLF)    . 
	--          The faces of the set theLF and theFace  must 
        --          share the edge theEdge  	
    	returns Boolean from Standard;  
	 
    IsInternalFace(myclass; 
    	    	theFace  :Face  from TopoDS; 
    	    	theSolid :Solid from TopoDS; 
		theMEF   :IndexedDataMapOfShapeListOfShape from TopTools;
    	    	theTol   :Real from Standard;       
    	    	theContext:out Context from IntTools)  
    	---Purpose: Returns True if the face theFace is inside the  
	--          solid theSolid. 
	--          theMEF - Map Edge/Faces for theSolid           	 
	--          theTol - value of precision of computation   
        --          theContext- cahed geometrical tools   
    	returns Boolean from Standard; 
    	
    
    GetFaceOff(myclass;  
    	    	theEdge    :Edge  from TopoDS;  
		theFace    :Face  from TopoDS; 
		theLCEF    :ListOfCoupleOfShape from NMTTools; 
		theFaceOff :out Face  from TopoDS); 
     	---Purpose:  For the face theFace and its edge theEdge 
        --           finds the face suitable to produce shell. 
	--           theLCEF - set of faces to search. All faces 
	--           from theLCEF must share edge theEdge 
	 
    GetEdgeOnFace (myclass;  
    	    	theEdge    :Edge  from TopoDS;  
		theFace    :Face  from TopoDS;  
		theEdgeOnF :out Edge  from TopoDS)  
	---Purpose: For the face theFace gets the edge theEdgeOnF 
        --          that is the same as theEdge 
        --          Returns True if such edge exists     	 
        --          Returns False if there is no such edge    	 
	returns Boolean from Standard; 
	 
    GetEdgeOff (myclass;  
    	    	theEdge    :Edge  from TopoDS;  
		theFace    :Face  from TopoDS;  
		theEdgeOff :out Edge  from TopoDS) 
    	---Purpose: Returns True if the face theFace contains 
	--          the edge theEdge but with opposite orientation. 
        --          If the method  returns True theEdgeOff is the 
        --          edge founded 	 
	returns Boolean from Standard; 

--fields
end Tools3D; 

