--  Copyright (C) 2007-2008  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--
-- File:	GEOMAlgo_GlueAnalyser.cdl
-- Created:	Wed Dec 15 11:03:03 2004
-- Author:	Peter KURNEV
--		<pkv@irinox>
--
class GlueAnalyser from GEOMAlgo 
    inherits Gluer from GEOMAlgo  
	---Purpose: 

uses 
    ShapeEnum from TopAbs, 
    ListOfShape from TopTools,
    ListOfCoupleOfShapes from GEOMAlgo

--raises

is
    Create   
    	returns GlueAnalyser from GEOMAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_GlueAnalyser();"

    Perform(me:out) 
	is redefined; 
	 
    HasSolidsToGlue(me)   
        returns Boolean from Standard;  
     
    SolidsToGlue(me) 
    	returns ListOfCoupleOfShapes from GEOMAlgo; 
    ---C++:return const &  
     
    HasSolidsAlone(me)   
        returns Boolean from Standard; 
     
    SolidsAlone(me) 
    	returns ListOfShape from TopTools; 
    ---C++:return const &   
     
    DetectVertices(me:out) 
	is protected;  
     
    DetectEdges(me:out) 
	is protected; 
     
    DetectFaces(me:out) 
	is protected;
     
    DetectShapes(me:out; 
    	    aType:ShapeEnum from TopAbs) 
    	is protected;        

    DetectSolids (me:out) 
    	is protected; 
	
    
     
fields  
    mySolidsToGlue   : ListOfCoupleOfShapes from GEOMAlgo is protected; 
    mySolidsAlone    : ListOfShape from TopTools is protected; 
    
end GlueAnalyser;
